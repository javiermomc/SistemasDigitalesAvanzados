----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:38:43 09/11/2019 
-- Design Name: 
-- Module Name:    Ones_Counter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Ones_Counter is
	 Generic ( n: integer:=7);
    Port ( A : in  STD_LOGIC_VECTOR (7 downto 0);
           SEG : out  STD_LOGIC_VECTOR (7 downto 0);
           ANODE : out  STD_LOGIC_VECTOR (3 downto 0));
end Ones_Counter;

architecture Behavioral of Ones_Counter is

signal BIN: STD_LOGIC_VECTOR(3 downto 0);

begin
	ANODE <= "0001";
	
	BIN <= ("000"&A(0))+("000"&A(1))+("000"&A(2))+("000"&A(3))+("000"&A(4))+("000"&A(5))+("000"&A(6))+("000"&A(7));
	with BIN select
      Seg <= x"C0" when x"0",
             x"F9" when x"1",
				 x"A4" when x"2",
				 x"B0" when x"3",
				 x"99" when x"4",
				 x"92" when x"5",
				 x"82" when x"6",
				 x"F8" when x"7",
				 x"80" when x"8",
				 x"90" when x"9",
				 x"88" when x"A",
				 x"83" when x"B",
				 x"C6" when x"C",
				 x"A1" when x"D",
				 x"86" when x"E",
				 x"8E" when x"F",
             x"7F" when others;
	
end Behavioral;

